module vga_controller (
  input logic clk,
  input logic rst,
  input logic perceptron_output,
  output logic[3:0] red,
  output logic[3:0] green,
  output logic[3:0] blue
);

endmodule
