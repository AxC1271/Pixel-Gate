module memory_interface (
  input logic clk,
  input logic rst,
  output logic[7:0] pixel_data,
  output logic valid
);

  
endmodule
