module graphics_driver (
  input logic clk,
  input logic rst,
  output logic[3:0] red,
  output logic[3:0] green,
  output logic[3:0] blue
);

end module;
